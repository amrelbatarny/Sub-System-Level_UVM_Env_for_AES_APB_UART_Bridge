package bridge_pkg;
    import uvm_pkg::*;
    import shared_pkg::*;
    `include "uvm_macros.svh"
    `include "agent_typedefs.svh"

    // Sequence Items
    `include "sequence_items/APB_sequence_item_base.svh"
    `include "sequence_items/APB_sequence_item_1.svh"
    `include "sequence_items/APB_sequence_item_2.svh"
    `include "sequence_items/APB_controller_sequence_item.svh"
    `include "sequence_items/AES_sequence_item.svh"
    `include "sequence_items/SYSCTRL_sequence_item.svh"
    
    // Sequencers
    `include "sequencers/APB_sequencer.svh"
    `include "sequencers/AES_sequencer.svh"
    `include "sequencers/SYSCTRL_sequencer.svh"

    // Sequencer Pool (Singleton Class)
    `include "sequencer_pool.svh"

    // Configuration Objects
    `include "env_config.svh"
    `include "agent_config.svh"

    // Monitors
    `include "monitors/APB_monitor_base.svh"
    `include "monitors/APB_monitor.svh"
    `include "monitors/APB_controller_monitor.svh"
    `include "monitors/AES_monitor.svh"
    `include "monitors/SYSCTRL_monitor.svh"

    // Drivers
    `include "drivers/APB_driver_base.svh"
    `include "drivers/APB_driver_1.svh"
    `include "drivers/APB_driver_2.svh"
    `include "drivers/SYSCTRL_driver.svh"
    `include "drivers/dummy_driver.svh"
    
    // Agent (Generic/Parameterized)
    `include "agent.svh"
    
    // Scoreboards
    `include "scoreboards/scoreboard_base.svh"
    `include "scoreboards/APB_scoreboard.svh"
    `include "scoreboards/APB_controller_scoreboard.svh"
    `include "scoreboards/AES_scoreboard.svh"

    // Environment
    `include "env.svh"
    
    // Base Sequences
    `include "virtual_sequence/virtual_sequence_base.svh"
    `include "reactive_sequences/APB_sequence_base.svh"

    // Reactive Sequences
    `include "reactive_sequences/APB_reactive_sequence_1.svh"
    `include "reactive_sequences/APB_reactive_sequence_2.svh"
    `include "virtual_sequence/virtual_sequence.svh"
    
    // Tests    
    `include "bridge_test_base.svh"
    
endpackage : bridge_pkg
